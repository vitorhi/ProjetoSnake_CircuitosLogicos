-------------------------------------------------------------------------------
--
-- Title       : 
-- Design      : Snake
-- Author      : Wang
--
-------------------------------------------------------------------------------
--
-- Description : 	Map/mask for the memory contents (VGA screen)
--					
--				Given the type of object in main memory , to output the corresponding map
-------------------------------------------------------------------------------


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.ALL;
use work.snake_package.all;
use work.vga_package.all;


entity all_maps is 
port	(
	my_code				: in code;						--data code in memory
	match_map			: out template_map 					--sketch to screen
	);
end all_maps;



architecture arch of all_maps is



signal blank_map_s:  template_map :=
("00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000");


signal body_map_s:  template_map :=
("00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
);

signal head_up_map_s:  template_map :=
("00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000011000000000000000"
,"00000000000000011000000000000000"
,"00000000000000111100000000000000"
,"00000000000000111100000000000000"
,"00000000000001111110000000000000"
,"00000000000001111110000000000000"
,"00000000000011111111000000000000"
,"00000000000011111111000000000000"
,"00000000000111111111100000000000"
,"00000000000111111111100000000000"
,"00000000001111111111110000000000"
,"00000000001111111111110000000000"
,"00000000011111111111111000000000"
,"00000000011111111111111000000000"
,"00000000111111111111111100000000"
,"00000000111111111111111100000000"
,"00000001111111111111111110000000"
,"00000001111111111111111110000000"
,"00000011111111111111111111000000"
,"00000011111111111111111111000000"
,"00000111111111111111111111100000"
,"00000111111111111111111111100000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000");

signal head_down_map_s:  template_map :=
("00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00000111111111111111111111100000"
,"00000111111111111111111111100000"
,"00000011111111111111111111000000"
,"00000011111111111111111111000000"
,"00000001111111111111111110000000"
,"00000001111111111111111110000000"
,"00000000111111111111111100000000"
,"00000000111111111111111100000000"
,"00000000011111111111111000000000"
,"00000000011111111111111000000000"
,"00000000001111111111110000000000"
,"00000000001111111111110000000000"
,"00000000000111111111100000000000"
,"00000000000111111111100000000000"
,"00000000000011111111000000000000"
,"00000000000011111111000000000000"
,"00000000000001111110000000000000"
,"00000000000001111110000000000000"
,"00000000000000111100000000000000"
,"00000000000000111100000000000000"
,"00000000000000011000000000000000"
,"00000000000000011000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000");

-- looks inverted due to the LSB/MSB placement
signal head_right_map_s:  template_map :=
("00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000110000"
,"00000000000000000000000011110000"
,"00000000000000000000001111110000"
,"00000000000000000000111111110000"
,"00000000000000000011111111110000"
,"00000000000000001111111111110000"
,"00000000000000111111111111110000"
,"00000000000011111111111111110000"
,"00000000001111111111111111110000"
,"00000000111111111111111111110000"
,"00000011111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00000011111111111111111111110000"
,"00000000111111111111111111110000"
,"00000000001111111111111111110000"
,"00000000000011111111111111110000"
,"00000000000000111111111111110000"
,"00000000000000001111111111110000"
,"00000000000000000011111111110000"
,"00000000000000000000111111110000"
,"00000000000000000000001111110000"
,"00000000000000000000000011110000"
,"00000000000000000000000000110000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000");


-- looks inverted due to the LSB/MSB placement
signal head_left_map_s:  template_map :=
("00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00001100000000000000000000000000"
,"00001111000000000000000000000000"
,"00001111110000000000000000000000"
,"00001111111100000000000000000000"
,"00001111111111000000000000000000"
,"00001111111111110000000000000000"
,"00001111111111111100000000000000"
,"00001111111111111111000000000000"
,"00001111111111111111110000000000"
,"00001111111111111111111100000000"
,"00001111111111111111111111000000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00001111111111111111111111000000"
,"00001111111111111111111100000000"
,"00001111111111111111110000000000"
,"00001111111111111111000000000000"
,"00001111111111111100000000000000"
,"00001111111111110000000000000000"
,"00001111111111000000000000000000"
,"00001111111100000000000000000000"
,"00001111110000000000000000000000"
,"00001111000000000000000000000000"
,"00001100000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000");

signal food_map_s:  template_map :=
("00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000111000000000111100000000"
,"00000011111110000001111111000000"
,"00000111111111000011111111100000"
,"00000111111111000011111111100000"
,"00001111111111000011111111110000"
,"00001111111111100111111111110000"
,"00000011111111111111111111000000"
,"00000000111111111111111100000000"
,"00000001111111111111111110000000"
,"00000001111111111111111110000000"
,"00000001111111111111111110000000"
,"00000011111111111111111111000000"
,"00000111111111111111111111100000"
,"00001111111111111111111111110000"
,"00001111111111111111111111110000"
,"00000011111111111111111111000000"
,"00000011111111111111111111000000"
,"00000011111111111111111111000000"
,"00000001111111111111111110000000"
,"00000000111111111111111100000000"
,"00000000011111111111111000000000"
,"00000000111111111111111100000000"
,"00000000001111100111110000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000"
,"00000000000000000000000000000000");


begin

	match_map <= 	blank_map_s when (my_code = BLANK) else
				food_map_s when (my_code = FOOD) else					
				body_map_s when (my_code = S_BODY) else 				
				head_up_map_s when (my_code = HEAD_UP) else	
				head_down_map_s when (my_code = HEAD_DOWN) else	
				head_right_map_s when (my_code = HEAD_RIGHT) else	
				head_left_map_s when (my_code = HEAD_LEFT);		
	
end arch;
